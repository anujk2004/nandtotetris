`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:15:07 05/14/2025 
// Design Name: 
// Module Name:    or16 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module or16(a,b,c
    );
input [0:8] a;
input [0:8] b;
output [0:8]c;

assign c= a||b;

endmodule
